module sdc_controller(clk, led, switch[7:0],  )
	reg [2:0] ch_sel;
	